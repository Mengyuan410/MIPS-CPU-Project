module pipe_alu (
    input logic clk,
    input logic waitrequest,
    input logic AluRegEn,
    input logic[3:0] AluControl,
    input logic[31:0] AluSrcIn1,
    input logic[31:0] AluSrcIn2,
    input logic AluSrc2Sel,
    input logic [31:0] Instruction,
    output logic[63:0] ALU // output can be even bigger
);
    logic [31:0] Immediate;
    logic [5:0] Opcode;
    logic [5:0] Funccode;
    logic [31:0] SignedImmediate, UnsignedImmediate;
    logic signed [31:0] SignedAluSrc1;
    logic signed [31:0] SignedAluSrc2;
    logic [31:0] AluSrc1, AluSrc2;
    logic [63:0] Result;

    assign Opcode = Instruction[31:26];
    assign Funccode = Instruction[5:0];
    assign UnsignedImmediate = Instruction[15:0];
    assign SignedImmediate =  {{16{Instruction[15]}}, (Instruction[15:0])};
    assign Immediate = ((Opcode[5]==1) || (Opcode == 6'b001001)|| (Opcode == 6'b001010) || (Opcode == 6'b001011)) ? SignedImmediate : UnsignedImmediate; //immediate is signed for load store
    assign AluSrc2= (AluSrc2Sel)? Immediate : AluSrcIn2;   
    assign AluSrc1 = (Opcode == 0 && Funccode[5:2] ==0)? AluSrcIn2 : AluSrcIn1; 
    assign SignedAluSrc1 = AluSrc1;
    assign SignedAluSrc2 = AluSrc2;

    always @(*) begin
        if (AluControl == 4'b0000) begin
            Result = AluSrc1 & AluSrc2; // AND 
        end
        
        else if (AluControl == 4'b0001) begin
            Result = AluSrc1 | AluSrc2; // OR and ORI
        end
        
        else if (AluControl == 4'b0010) begin
            Result = AluSrc1 + AluSrc2; //for the add and since the operation codes are the same for LW and SW
        end
        
        else if(AluControl == 4'b0011 )begin // SLL SLLV
            if(AluSrc2Sel == 0)begin
                //SLLV
                Result = AluSrc2 << AluSrc1;
            end
            else begin
                //SLL
                Result = AluSrc1 << AluSrc2[10:6];
            end

        end
        else if(AluControl == 4'b0100) begin // SLTU
            Result = (AluSrc1 < AluSrc2);
        end
        else if(AluControl == 4'b0101) begin // SRA SRAV
            if(AluSrc2Sel == 0)begin
                //SRAV
                Result[31:0] = SignedAluSrc2 >>> SignedAluSrc1;
            end
            else begin
                //SRA
                Result = SignedAluSrc1 >>> SignedAluSrc2[10:6];
            end
        end
        else if(AluControl == 4'b0110) begin // SUBU
            Result = AluSrc1 - AluSrc2;
        end
        else if(AluControl == 4'b0111) begin // SLT SLTI
            Result = (SignedAluSrc1 < SignedAluSrc2);
        end
        else if(AluControl == 4'b1000) begin // divide signed
            Result[31:0] = SignedAluSrc1 / SignedAluSrc2;
            Result[63:32] = SignedAluSrc1 % SignedAluSrc2;
        end
        else if(AluControl == 4'b1001) begin // divide unsigned
            Result[31:0] = AluSrc1 / AluSrc2;
            Result[63:32] = AluSrc1 % AluSrc2;
        end
        
        else if(AluControl == 4'b1010) begin // multiply signed
            Result = SignedAluSrc1 * SignedAluSrc2;
        end
        
        else if(AluControl == 4'b1011) begin // multiply unsigned
            Result = AluSrc1 * AluSrc2;
        end
        
        else if(AluControl == 4'b1100) begin // shift right logical
            if(AluSrc2Sel == 0)begin //SRLV
                Result = AluSrc2 >> AluSrc1;
            end
            else begin //SRL
                Result = AluSrc1 >> AluSrc2[10:6];
            end
        end

        else if(AluControl == 4'b1101) begin // XOR
            Result = AluSrc1 ^ AluSrc2; 
        end
        else if(AluControl == 4'b1110) begin // LUI
            Result = AluSrc2 << 16; 
        end
        else if(AluControl == 4'b1111) begin // do nothing
            Result = 32'hxxxxxxxx;
        end
    end


    always_ff @(posedge clk) begin
        if (AluRegEn==1 && waitrequest == 0)begin
            ALU <= Result;
        end
    end

endmodule

